// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Mon Sep 27 11:57:43 2021
//
// Verilog Description of module distance_ram
//

module distance_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(8[8:20])
    input [7:0]WrAddress;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(10[22:31])
    input [7:0]RdAddress;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(11[22:31])
    input [63:0]Data;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(12[23:27])
    input WE;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(13[16:18])
    input RdClock;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(14[16:23])
    input RdClockEn;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(15[16:25])
    input Reset;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(16[16:21])
    input WrClock;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(17[16:23])
    input WrClockEn;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(18[16:25])
    output [63:0]Q;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(19[24:25])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c252/c25x_21092711_encoder/c25x_fpga_ip/distance_ram/distance_ram.v(17[16:23])
    
    wire scuba_vlo, VCC_net;
    
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    PDPW16KD distance_ram_0_1_0 (.DI0(Data[36]), .DI1(Data[37]), .DI2(Data[38]), 
            .DI3(Data[39]), .DI4(Data[40]), .DI5(Data[41]), .DI6(Data[42]), 
            .DI7(Data[43]), .DI8(Data[44]), .DI9(Data[45]), .DI10(Data[46]), 
            .DI11(Data[47]), .DI12(Data[48]), .DI13(Data[49]), .DI14(Data[50]), 
            .DI15(Data[51]), .DI16(Data[52]), .DI17(Data[53]), .DI18(Data[54]), 
            .DI19(Data[55]), .DI20(Data[56]), .DI21(Data[57]), .DI22(Data[58]), 
            .DI23(Data[59]), .DI24(Data[60]), .DI25(Data[61]), .DI26(Data[62]), 
            .DI27(Data[63]), .DI28(scuba_vlo), .DI29(scuba_vlo), .DI30(scuba_vlo), 
            .DI31(scuba_vlo), .DI32(scuba_vlo), .DI33(scuba_vlo), .DI34(scuba_vlo), 
            .DI35(scuba_vlo), .ADW0(WrAddress[0]), .ADW1(WrAddress[1]), 
            .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), .ADW4(WrAddress[4]), 
            .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), .ADW7(WrAddress[7]), 
            .ADW8(scuba_vlo), .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), 
            .BE3(VCC_net), .CEW(WrClockEn), .CLKW(WrClock), .CSW0(WE), 
            .CSW1(scuba_vlo), .CSW2(scuba_vlo), .ADR0(scuba_vlo), .ADR1(scuba_vlo), 
            .ADR2(scuba_vlo), .ADR3(scuba_vlo), .ADR4(scuba_vlo), .ADR5(RdAddress[0]), 
            .ADR6(RdAddress[1]), .ADR7(RdAddress[2]), .ADR8(RdAddress[3]), 
            .ADR9(RdAddress[4]), .ADR10(RdAddress[5]), .ADR11(RdAddress[6]), 
            .ADR12(RdAddress[7]), .ADR13(scuba_vlo), .CER(RdClockEn), 
            .OCER(RdClockEn), .CLKR(RdClock), .CSR0(scuba_vlo), .CSR1(scuba_vlo), 
            .CSR2(scuba_vlo), .RST(Reset), .DO0(Q[54]), .DO1(Q[55]), 
            .DO2(Q[56]), .DO3(Q[57]), .DO4(Q[58]), .DO5(Q[59]), .DO6(Q[60]), 
            .DO7(Q[61]), .DO8(Q[62]), .DO9(Q[63]), .DO18(Q[36]), .DO19(Q[37]), 
            .DO20(Q[38]), .DO21(Q[39]), .DO22(Q[40]), .DO23(Q[41]), 
            .DO24(Q[42]), .DO25(Q[43]), .DO26(Q[44]), .DO27(Q[45]), 
            .DO28(Q[46]), .DO29(Q[47]), .DO30(Q[48]), .DO31(Q[49]), 
            .DO32(Q[50]), .DO33(Q[51]), .DO34(Q[52]), .DO35(Q[53])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_1_0.DATA_WIDTH_W = 36;
    defparam distance_ram_0_1_0.DATA_WIDTH_R = 36;
    defparam distance_ram_0_1_0.GSR = "ENABLED";
    defparam distance_ram_0_1_0.REGMODE = "NOREG";
    defparam distance_ram_0_1_0.RESETMODE = "ASYNC";
    defparam distance_ram_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_1_0.CSDECODE_W = "0b001";
    defparam distance_ram_0_1_0.CSDECODE_R = "0b000";
    defparam distance_ram_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_0.INIT_DATA = "STATIC";
    PDPW16KD distance_ram_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .DI18(Data[18]), 
            .DI19(Data[19]), .DI20(Data[20]), .DI21(Data[21]), .DI22(Data[22]), 
            .DI23(Data[23]), .DI24(Data[24]), .DI25(Data[25]), .DI26(Data[26]), 
            .DI27(Data[27]), .DI28(Data[28]), .DI29(Data[29]), .DI30(Data[30]), 
            .DI31(Data[31]), .DI32(Data[32]), .DI33(Data[33]), .DI34(Data[34]), 
            .DI35(Data[35]), .ADW0(WrAddress[0]), .ADW1(WrAddress[1]), 
            .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), .ADW4(WrAddress[4]), 
            .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), .ADW7(WrAddress[7]), 
            .ADW8(scuba_vlo), .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), 
            .BE3(VCC_net), .CEW(WrClockEn), .CLKW(WrClock), .CSW0(WE), 
            .CSW1(scuba_vlo), .CSW2(scuba_vlo), .ADR0(scuba_vlo), .ADR1(scuba_vlo), 
            .ADR2(scuba_vlo), .ADR3(scuba_vlo), .ADR4(scuba_vlo), .ADR5(RdAddress[0]), 
            .ADR6(RdAddress[1]), .ADR7(RdAddress[2]), .ADR8(RdAddress[3]), 
            .ADR9(RdAddress[4]), .ADR10(RdAddress[5]), .ADR11(RdAddress[6]), 
            .ADR12(RdAddress[7]), .ADR13(scuba_vlo), .CER(RdClockEn), 
            .OCER(RdClockEn), .CLKR(RdClock), .CSR0(scuba_vlo), .CSR1(scuba_vlo), 
            .CSR2(scuba_vlo), .RST(Reset), .DO0(Q[18]), .DO1(Q[19]), 
            .DO2(Q[20]), .DO3(Q[21]), .DO4(Q[22]), .DO5(Q[23]), .DO6(Q[24]), 
            .DO7(Q[25]), .DO8(Q[26]), .DO9(Q[27]), .DO10(Q[28]), .DO11(Q[29]), 
            .DO12(Q[30]), .DO13(Q[31]), .DO14(Q[32]), .DO15(Q[33]), 
            .DO16(Q[34]), .DO17(Q[35]), .DO18(Q[0]), .DO19(Q[1]), .DO20(Q[2]), 
            .DO21(Q[3]), .DO22(Q[4]), .DO23(Q[5]), .DO24(Q[6]), .DO25(Q[7]), 
            .DO26(Q[8]), .DO27(Q[9]), .DO28(Q[10]), .DO29(Q[11]), .DO30(Q[12]), 
            .DO31(Q[13]), .DO32(Q[14]), .DO33(Q[15]), .DO34(Q[16]), 
            .DO35(Q[17])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_0_1.DATA_WIDTH_W = 36;
    defparam distance_ram_0_0_1.DATA_WIDTH_R = 36;
    defparam distance_ram_0_0_1.GSR = "ENABLED";
    defparam distance_ram_0_0_1.REGMODE = "NOREG";
    defparam distance_ram_0_0_1.RESETMODE = "ASYNC";
    defparam distance_ram_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_0_1.CSDECODE_W = "0b001";
    defparam distance_ram_0_0_1.CSDECODE_R = "0b000";
    defparam distance_ram_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_1.INIT_DATA = "STATIC";
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VHI i157 (.Z(VCC_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

