// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Sat Mar 29 16:30:09 2025
//
// Verilog Description of module cache_opto_ram
//

module cache_opto_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(8[8:22])
    input [7:0]WrAddress;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(10[22:31])
    input [7:0]RdAddress;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(11[22:31])
    input [15:0]Data;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(12[23:27])
    input WE;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(13[16:18])
    input RdClock;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(14[16:23])
    input RdClockEn;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(15[16:25])
    input Reset;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(16[16:21])
    input WrClock;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(17[16:23])
    input WrClockEn;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(18[16:25])
    output [15:0]Q;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(19[24:25])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200/h100/h100_fpga/c25x_fpga_ip/cache_opto_ram/cache_opto_ram.v(17[16:23])
    
    wire scuba_vlo, VCC_net;
    
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    DP16KD cache_opto_ram_0_0_0_0 (.DIA0(Data[0]), .DIA1(Data[1]), .DIA2(Data[2]), 
           .DIA3(Data[3]), .DIA4(Data[4]), .DIA5(Data[5]), .DIA6(Data[6]), 
           .DIA7(Data[7]), .DIA8(Data[8]), .DIA9(Data[9]), .DIA10(Data[10]), 
           .DIA11(Data[11]), .DIA12(Data[12]), .DIA13(Data[13]), .DIA14(Data[14]), 
           .DIA15(Data[15]), .DIA16(scuba_vlo), .DIA17(scuba_vlo), .ADA0(VCC_net), 
           .ADA1(VCC_net), .ADA2(scuba_vlo), .ADA3(scuba_vlo), .ADA4(WrAddress[0]), 
           .ADA5(WrAddress[1]), .ADA6(WrAddress[2]), .ADA7(WrAddress[3]), 
           .ADA8(WrAddress[4]), .ADA9(WrAddress[5]), .ADA10(WrAddress[6]), 
           .ADA11(WrAddress[7]), .ADA12(scuba_vlo), .ADA13(scuba_vlo), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset), 
           .DIB0(scuba_vlo), .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), 
           .DIB4(scuba_vlo), .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), 
           .DIB8(scuba_vlo), .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), 
           .DIB12(scuba_vlo), .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), 
           .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), 
           .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(RdAddress[0]), .ADB5(RdAddress[1]), 
           .ADB6(RdAddress[2]), .ADB7(RdAddress[3]), .ADB8(RdAddress[4]), 
           .ADB9(RdAddress[5]), .ADB10(RdAddress[6]), .ADB11(RdAddress[7]), 
           .ADB12(scuba_vlo), .ADB13(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), 
           .CLKB(RdClock), .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), 
           .CSB2(scuba_vlo), .RSTB(Reset), .DOB0(Q[0]), .DOB1(Q[1]), 
           .DOB2(Q[2]), .DOB3(Q[3]), .DOB4(Q[4]), .DOB5(Q[5]), .DOB6(Q[6]), 
           .DOB7(Q[7]), .DOB8(Q[8]), .DOB9(Q[9]), .DOB10(Q[10]), .DOB11(Q[11]), 
           .DOB12(Q[12]), .DOB13(Q[13]), .DOB14(Q[14]), .DOB15(Q[15])) /* synthesis MEM_LPC_FILE="cache_opto_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam cache_opto_ram_0_0_0_0.DATA_WIDTH_A = 18;
    defparam cache_opto_ram_0_0_0_0.DATA_WIDTH_B = 18;
    defparam cache_opto_ram_0_0_0_0.REGMODE_A = "NOREG";
    defparam cache_opto_ram_0_0_0_0.REGMODE_B = "NOREG";
    defparam cache_opto_ram_0_0_0_0.RESETMODE = "ASYNC";
    defparam cache_opto_ram_0_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam cache_opto_ram_0_0_0_0.WRITEMODE_A = "NORMAL";
    defparam cache_opto_ram_0_0_0_0.WRITEMODE_B = "NORMAL";
    defparam cache_opto_ram_0_0_0_0.CSDECODE_A = "0b000";
    defparam cache_opto_ram_0_0_0_0.CSDECODE_B = "0b000";
    defparam cache_opto_ram_0_0_0_0.GSR = "ENABLED";
    defparam cache_opto_ram_0_0_0_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam cache_opto_ram_0_0_0_0.INIT_DATA = "STATIC";
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VHI i60 (.Z(VCC_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

