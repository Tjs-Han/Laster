// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Wed Dec 14 10:10:16 2022
//
// Verilog Description of module tcp_recv_ram
//

module tcp_recv_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(8[8:20])
    input [11:0]WrAddress;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(10[23:32])
    input [11:0]RdAddress;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(11[23:32])
    input [7:0]Data;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(12[22:26])
    input WE;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(13[16:18])
    input RdClock;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(14[16:23])
    input RdClockEn;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(15[16:25])
    input Reset;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(16[16:21])
    input WrClock;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(17[16:23])
    input WrClockEn;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(18[16:25])
    output [7:0]Q;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(19[23:24])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // c:/users/guoxiang/desktop/fpga/c200/program_formal/c200/haikang/c200_fpga_gp22_22090813/c200_fpga/tcp_recv_ram/tcp_recv_ram.v(17[16:23])
    
    wire GND_net, VCC_net;
    
    DP16KD tcp_recv_ram_0_0_1 (.DIA0(Data[0]), .DIA1(Data[1]), .DIA2(Data[2]), 
           .DIA3(Data[3]), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
           .DIA7(GND_net), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(WrAddress[0]), .ADA3(WrAddress[1]), .ADA4(WrAddress[2]), 
           .ADA5(WrAddress[3]), .ADA6(WrAddress[4]), .ADA7(WrAddress[5]), 
           .ADA8(WrAddress[6]), .ADA9(WrAddress[7]), .ADA10(WrAddress[8]), 
           .ADA11(WrAddress[9]), .ADA12(WrAddress[10]), .ADA13(WrAddress[11]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(RdAddress[0]), .ADB3(RdAddress[1]), .ADB4(RdAddress[2]), 
           .ADB5(RdAddress[3]), .ADB6(RdAddress[4]), .ADB7(RdAddress[5]), 
           .ADB8(RdAddress[6]), .ADB9(RdAddress[7]), .ADB10(RdAddress[8]), 
           .ADB11(RdAddress[9]), .ADB12(RdAddress[10]), .ADB13(RdAddress[11]), 
           .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), 
           .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), 
           .DOB0(Q[0]), .DOB1(Q[1]), .DOB2(Q[2]), .DOB3(Q[3])) /* synthesis MEM_LPC_FILE="tcp_recv_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam tcp_recv_ram_0_0_1.DATA_WIDTH_A = 4;
    defparam tcp_recv_ram_0_0_1.DATA_WIDTH_B = 4;
    defparam tcp_recv_ram_0_0_1.REGMODE_A = "OUTREG";
    defparam tcp_recv_ram_0_0_1.REGMODE_B = "OUTREG";
    defparam tcp_recv_ram_0_0_1.RESETMODE = "SYNC";
    defparam tcp_recv_ram_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam tcp_recv_ram_0_0_1.WRITEMODE_A = "NORMAL";
    defparam tcp_recv_ram_0_0_1.WRITEMODE_B = "NORMAL";
    defparam tcp_recv_ram_0_0_1.CSDECODE_A = "0b000";
    defparam tcp_recv_ram_0_0_1.CSDECODE_B = "0b000";
    defparam tcp_recv_ram_0_0_1.GSR = "ENABLED";
    defparam tcp_recv_ram_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_0_1.INIT_DATA = "STATIC";
    DP16KD tcp_recv_ram_0_1_0 (.DIA0(Data[4]), .DIA1(Data[5]), .DIA2(Data[6]), 
           .DIA3(Data[7]), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
           .DIA7(GND_net), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(WrAddress[0]), .ADA3(WrAddress[1]), .ADA4(WrAddress[2]), 
           .ADA5(WrAddress[3]), .ADA6(WrAddress[4]), .ADA7(WrAddress[5]), 
           .ADA8(WrAddress[6]), .ADA9(WrAddress[7]), .ADA10(WrAddress[8]), 
           .ADA11(WrAddress[9]), .ADA12(WrAddress[10]), .ADA13(WrAddress[11]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(RdAddress[0]), .ADB3(RdAddress[1]), .ADB4(RdAddress[2]), 
           .ADB5(RdAddress[3]), .ADB6(RdAddress[4]), .ADB7(RdAddress[5]), 
           .ADB8(RdAddress[6]), .ADB9(RdAddress[7]), .ADB10(RdAddress[8]), 
           .ADB11(RdAddress[9]), .ADB12(RdAddress[10]), .ADB13(RdAddress[11]), 
           .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), 
           .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), 
           .DOB0(Q[4]), .DOB1(Q[5]), .DOB2(Q[6]), .DOB3(Q[7])) /* synthesis MEM_LPC_FILE="tcp_recv_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam tcp_recv_ram_0_1_0.DATA_WIDTH_A = 4;
    defparam tcp_recv_ram_0_1_0.DATA_WIDTH_B = 4;
    defparam tcp_recv_ram_0_1_0.REGMODE_A = "OUTREG";
    defparam tcp_recv_ram_0_1_0.REGMODE_B = "OUTREG";
    defparam tcp_recv_ram_0_1_0.RESETMODE = "SYNC";
    defparam tcp_recv_ram_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam tcp_recv_ram_0_1_0.WRITEMODE_A = "NORMAL";
    defparam tcp_recv_ram_0_1_0.WRITEMODE_B = "NORMAL";
    defparam tcp_recv_ram_0_1_0.CSDECODE_A = "0b000";
    defparam tcp_recv_ram_0_1_0.CSDECODE_B = "0b000";
    defparam tcp_recv_ram_0_1_0.GSR = "ENABLED";
    defparam tcp_recv_ram_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tcp_recv_ram_0_1_0.INIT_DATA = "STATIC";
    VHI i13 (.Z(VCC_net));
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i4 (.Z(GND_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

