// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Tue Jun 15 14:32:02 2021
//
// Verilog Description of module eth_send_ram
//

module eth_send_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(8[8:20])
    input [10:0]WrAddress;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(10[23:32])
    input [10:0]RdAddress;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(11[23:32])
    input [7:0]Data;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(12[22:26])
    input WE;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(13[16:18])
    input RdClock;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(14[16:23])
    input RdClockEn;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(15[16:25])
    input Reset;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(16[16:21])
    input WrClock;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(17[16:23])
    input WrClockEn;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(18[16:25])
    output [7:0]Q;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(19[23:24])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/eth_send_ram/eth_send_ram.v(17[16:23])
    
    wire scuba_vlo, VCC_net;
    
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    DP16KD eth_send_ram_0_0_0 (.DIA0(Data[0]), .DIA1(Data[1]), .DIA2(Data[2]), 
           .DIA3(Data[3]), .DIA4(Data[4]), .DIA5(Data[5]), .DIA6(Data[6]), 
           .DIA7(Data[7]), .DIA8(scuba_vlo), .DIA9(scuba_vlo), .DIA10(scuba_vlo), 
           .DIA11(scuba_vlo), .DIA12(scuba_vlo), .DIA13(scuba_vlo), .DIA14(scuba_vlo), 
           .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), .ADA0(scuba_vlo), 
           .ADA1(scuba_vlo), .ADA2(scuba_vlo), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset), 
           .DIB0(scuba_vlo), .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), 
           .DIB4(scuba_vlo), .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), 
           .DIB8(scuba_vlo), .DIB9(scuba_vlo), .DIB10(scuba_vlo), .DIB11(scuba_vlo), 
           .DIB12(scuba_vlo), .DIB13(scuba_vlo), .DIB14(scuba_vlo), .DIB15(scuba_vlo), 
           .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vlo), .ADB1(scuba_vlo), 
           .ADB2(scuba_vlo), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), 
           .ADB5(RdAddress[2]), .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), 
           .ADB8(RdAddress[5]), .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), 
           .ADB11(RdAddress[8]), .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), 
           .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
           .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), .RSTB(Reset), 
           .DOB0(Q[0]), .DOB1(Q[1]), .DOB2(Q[2]), .DOB3(Q[3]), .DOB4(Q[4]), 
           .DOB5(Q[5]), .DOB6(Q[6]), .DOB7(Q[7])) /* synthesis MEM_LPC_FILE="eth_send_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam eth_send_ram_0_0_0.DATA_WIDTH_A = 9;
    defparam eth_send_ram_0_0_0.DATA_WIDTH_B = 9;
    defparam eth_send_ram_0_0_0.REGMODE_A = "NOREG";
    defparam eth_send_ram_0_0_0.REGMODE_B = "NOREG";
    defparam eth_send_ram_0_0_0.RESETMODE = "ASYNC";
    defparam eth_send_ram_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam eth_send_ram_0_0_0.WRITEMODE_A = "NORMAL";
    defparam eth_send_ram_0_0_0.WRITEMODE_B = "NORMAL";
    defparam eth_send_ram_0_0_0.CSDECODE_A = "0b000";
    defparam eth_send_ram_0_0_0.CSDECODE_B = "0b000";
    defparam eth_send_ram_0_0_0.GSR = "ENABLED";
    defparam eth_send_ram_0_0_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam eth_send_ram_0_0_0.INIT_DATA = "STATIC";
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VHI i57 (.Z(VCC_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

