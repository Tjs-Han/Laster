// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Sun Jun 06 19:09:20 2021
//
// Verilog Description of module distance_ram
//

module distance_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(8[8:20])
    input [10:0]WrAddress;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(10[23:32])
    input [10:0]RdAddress;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(11[23:32])
    input [63:0]Data;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(12[23:27])
    input WE;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(13[16:18])
    input RdClock;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(14[16:23])
    input RdClockEn;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(15[16:25])
    input Reset;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(16[16:21])
    input WrClock;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(17[16:23])
    input WrClockEn;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(18[16:25])
    output [63:0]Q;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(19[24:25])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // d:/programs/fpga/c200_fpga/c200_fpga/distance_ram/distance_ram.v(17[16:23])
    
    wire GND_net, VCC_net;
    
    DP16KD distance_ram_0_0_7 (.DIA0(Data[0]), .DIA1(Data[1]), .DIA2(Data[2]), 
           .DIA3(Data[3]), .DIA4(Data[4]), .DIA5(Data[5]), .DIA6(Data[6]), 
           .DIA7(Data[7]), .DIA8(Data[8]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[0]), 
           .DOB1(Q[1]), .DOB2(Q[2]), .DOB3(Q[3]), .DOB4(Q[4]), .DOB5(Q[5]), 
           .DOB6(Q[6]), .DOB7(Q[7]), .DOB8(Q[8])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_0_7.DATA_WIDTH_A = 9;
    defparam distance_ram_0_0_7.DATA_WIDTH_B = 9;
    defparam distance_ram_0_0_7.REGMODE_A = "OUTREG";
    defparam distance_ram_0_0_7.REGMODE_B = "OUTREG";
    defparam distance_ram_0_0_7.RESETMODE = "SYNC";
    defparam distance_ram_0_0_7.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_0_7.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_0_7.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_0_7.CSDECODE_A = "0b000";
    defparam distance_ram_0_0_7.CSDECODE_B = "0b000";
    defparam distance_ram_0_0_7.GSR = "ENABLED";
    defparam distance_ram_0_0_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_0_7.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_7_0 (.DIA0(Data[63]), .DIA1(GND_net), .DIA2(GND_net), 
           .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
           .DIA7(GND_net), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[63])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_7_0.DATA_WIDTH_A = 9;
    defparam distance_ram_0_7_0.DATA_WIDTH_B = 9;
    defparam distance_ram_0_7_0.REGMODE_A = "OUTREG";
    defparam distance_ram_0_7_0.REGMODE_B = "OUTREG";
    defparam distance_ram_0_7_0.RESETMODE = "SYNC";
    defparam distance_ram_0_7_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_7_0.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_7_0.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_7_0.CSDECODE_A = "0b000";
    defparam distance_ram_0_7_0.CSDECODE_B = "0b000";
    defparam distance_ram_0_7_0.GSR = "ENABLED";
    defparam distance_ram_0_7_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_7_0.INIT_DATA = "STATIC";
    VHI i19 (.Z(VCC_net));
    DP16KD distance_ram_0_1_6 (.DIA0(Data[9]), .DIA1(Data[10]), .DIA2(Data[11]), 
           .DIA3(Data[12]), .DIA4(Data[13]), .DIA5(Data[14]), .DIA6(Data[15]), 
           .DIA7(Data[16]), .DIA8(Data[17]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[9]), 
           .DOB1(Q[10]), .DOB2(Q[11]), .DOB3(Q[12]), .DOB4(Q[13]), .DOB5(Q[14]), 
           .DOB6(Q[15]), .DOB7(Q[16]), .DOB8(Q[17])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_1_6.DATA_WIDTH_A = 9;
    defparam distance_ram_0_1_6.DATA_WIDTH_B = 9;
    defparam distance_ram_0_1_6.REGMODE_A = "OUTREG";
    defparam distance_ram_0_1_6.REGMODE_B = "OUTREG";
    defparam distance_ram_0_1_6.RESETMODE = "SYNC";
    defparam distance_ram_0_1_6.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_1_6.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_1_6.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_1_6.CSDECODE_A = "0b000";
    defparam distance_ram_0_1_6.CSDECODE_B = "0b000";
    defparam distance_ram_0_1_6.GSR = "ENABLED";
    defparam distance_ram_0_1_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_1_6.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_2_5 (.DIA0(Data[18]), .DIA1(Data[19]), .DIA2(Data[20]), 
           .DIA3(Data[21]), .DIA4(Data[22]), .DIA5(Data[23]), .DIA6(Data[24]), 
           .DIA7(Data[25]), .DIA8(Data[26]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[18]), 
           .DOB1(Q[19]), .DOB2(Q[20]), .DOB3(Q[21]), .DOB4(Q[22]), .DOB5(Q[23]), 
           .DOB6(Q[24]), .DOB7(Q[25]), .DOB8(Q[26])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_2_5.DATA_WIDTH_A = 9;
    defparam distance_ram_0_2_5.DATA_WIDTH_B = 9;
    defparam distance_ram_0_2_5.REGMODE_A = "OUTREG";
    defparam distance_ram_0_2_5.REGMODE_B = "OUTREG";
    defparam distance_ram_0_2_5.RESETMODE = "SYNC";
    defparam distance_ram_0_2_5.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_2_5.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_2_5.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_2_5.CSDECODE_A = "0b000";
    defparam distance_ram_0_2_5.CSDECODE_B = "0b000";
    defparam distance_ram_0_2_5.GSR = "ENABLED";
    defparam distance_ram_0_2_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_2_5.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_3_4 (.DIA0(Data[27]), .DIA1(Data[28]), .DIA2(Data[29]), 
           .DIA3(Data[30]), .DIA4(Data[31]), .DIA5(Data[32]), .DIA6(Data[33]), 
           .DIA7(Data[34]), .DIA8(Data[35]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[27]), 
           .DOB1(Q[28]), .DOB2(Q[29]), .DOB3(Q[30]), .DOB4(Q[31]), .DOB5(Q[32]), 
           .DOB6(Q[33]), .DOB7(Q[34]), .DOB8(Q[35])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_3_4.DATA_WIDTH_A = 9;
    defparam distance_ram_0_3_4.DATA_WIDTH_B = 9;
    defparam distance_ram_0_3_4.REGMODE_A = "OUTREG";
    defparam distance_ram_0_3_4.REGMODE_B = "OUTREG";
    defparam distance_ram_0_3_4.RESETMODE = "SYNC";
    defparam distance_ram_0_3_4.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_3_4.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_3_4.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_3_4.CSDECODE_A = "0b000";
    defparam distance_ram_0_3_4.CSDECODE_B = "0b000";
    defparam distance_ram_0_3_4.GSR = "ENABLED";
    defparam distance_ram_0_3_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_3_4.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_4_3 (.DIA0(Data[36]), .DIA1(Data[37]), .DIA2(Data[38]), 
           .DIA3(Data[39]), .DIA4(Data[40]), .DIA5(Data[41]), .DIA6(Data[42]), 
           .DIA7(Data[43]), .DIA8(Data[44]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[36]), 
           .DOB1(Q[37]), .DOB2(Q[38]), .DOB3(Q[39]), .DOB4(Q[40]), .DOB5(Q[41]), 
           .DOB6(Q[42]), .DOB7(Q[43]), .DOB8(Q[44])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_4_3.DATA_WIDTH_A = 9;
    defparam distance_ram_0_4_3.DATA_WIDTH_B = 9;
    defparam distance_ram_0_4_3.REGMODE_A = "OUTREG";
    defparam distance_ram_0_4_3.REGMODE_B = "OUTREG";
    defparam distance_ram_0_4_3.RESETMODE = "SYNC";
    defparam distance_ram_0_4_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_4_3.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_4_3.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_4_3.CSDECODE_A = "0b000";
    defparam distance_ram_0_4_3.CSDECODE_B = "0b000";
    defparam distance_ram_0_4_3.GSR = "ENABLED";
    defparam distance_ram_0_4_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_4_3.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_5_2 (.DIA0(Data[45]), .DIA1(Data[46]), .DIA2(Data[47]), 
           .DIA3(Data[48]), .DIA4(Data[49]), .DIA5(Data[50]), .DIA6(Data[51]), 
           .DIA7(Data[52]), .DIA8(Data[53]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[45]), 
           .DOB1(Q[46]), .DOB2(Q[47]), .DOB3(Q[48]), .DOB4(Q[49]), .DOB5(Q[50]), 
           .DOB6(Q[51]), .DOB7(Q[52]), .DOB8(Q[53])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_5_2.DATA_WIDTH_A = 9;
    defparam distance_ram_0_5_2.DATA_WIDTH_B = 9;
    defparam distance_ram_0_5_2.REGMODE_A = "OUTREG";
    defparam distance_ram_0_5_2.REGMODE_B = "OUTREG";
    defparam distance_ram_0_5_2.RESETMODE = "SYNC";
    defparam distance_ram_0_5_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_5_2.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_5_2.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_5_2.CSDECODE_A = "0b000";
    defparam distance_ram_0_5_2.CSDECODE_B = "0b000";
    defparam distance_ram_0_5_2.GSR = "ENABLED";
    defparam distance_ram_0_5_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_5_2.INIT_DATA = "STATIC";
    DP16KD distance_ram_0_6_1 (.DIA0(Data[54]), .DIA1(Data[55]), .DIA2(Data[56]), 
           .DIA3(Data[57]), .DIA4(Data[58]), .DIA5(Data[59]), .DIA6(Data[60]), 
           .DIA7(Data[61]), .DIA8(Data[62]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[54]), 
           .DOB1(Q[55]), .DOB2(Q[56]), .DOB3(Q[57]), .DOB4(Q[58]), .DOB5(Q[59]), 
           .DOB6(Q[60]), .DOB7(Q[61]), .DOB8(Q[62])) /* synthesis MEM_LPC_FILE="distance_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam distance_ram_0_6_1.DATA_WIDTH_A = 9;
    defparam distance_ram_0_6_1.DATA_WIDTH_B = 9;
    defparam distance_ram_0_6_1.REGMODE_A = "OUTREG";
    defparam distance_ram_0_6_1.REGMODE_B = "OUTREG";
    defparam distance_ram_0_6_1.RESETMODE = "SYNC";
    defparam distance_ram_0_6_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam distance_ram_0_6_1.WRITEMODE_A = "NORMAL";
    defparam distance_ram_0_6_1.WRITEMODE_B = "NORMAL";
    defparam distance_ram_0_6_1.CSDECODE_A = "0b000";
    defparam distance_ram_0_6_1.CSDECODE_B = "0b000";
    defparam distance_ram_0_6_1.GSR = "ENABLED";
    defparam distance_ram_0_6_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam distance_ram_0_6_1.INIT_DATA = "STATIC";
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i4 (.Z(GND_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

