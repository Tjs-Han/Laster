// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Sun Nov 28 13:20:35 2021
//
// Verilog Description of module tdc_data_ram
//

module tdc_data_ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, 
            Reset, WrClock, WrClockEn, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(8[8:20])
    input [10:0]WrAddress;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(10[23:32])
    input [10:0]RdAddress;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(11[23:32])
    input [15:0]Data;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(12[23:27])
    input WE;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(13[16:18])
    input RdClock;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(14[16:23])
    input RdClockEn;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(15[16:25])
    input Reset;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(16[16:21])
    input WrClock;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(17[16:23])
    input WrClockEn;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(18[16:25])
    output [15:0]Q;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(19[24:25])
    
    wire RdClock /* synthesis is_clock=1 */ ;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(14[16:23])
    wire WrClock /* synthesis is_clock=1 */ ;   // c:/users/guoxiang/desktop/c200/program_test/c200_fpga_gp22_20211128_temp/tdc_data/tdc_data_ram/tdc_data_ram.v(17[16:23])
    
    wire GND_net, VCC_net;
    
    DP16KD tdc_data_ram_0_0_1 (.DIA0(Data[0]), .DIA1(Data[1]), .DIA2(Data[2]), 
           .DIA3(Data[3]), .DIA4(Data[4]), .DIA5(Data[5]), .DIA6(Data[6]), 
           .DIA7(Data[7]), .DIA8(Data[8]), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[0]), 
           .DOB1(Q[1]), .DOB2(Q[2]), .DOB3(Q[3]), .DOB4(Q[4]), .DOB5(Q[5]), 
           .DOB6(Q[6]), .DOB7(Q[7]), .DOB8(Q[8])) /* synthesis MEM_LPC_FILE="tdc_data_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam tdc_data_ram_0_0_1.DATA_WIDTH_A = 9;
    defparam tdc_data_ram_0_0_1.DATA_WIDTH_B = 9;
    defparam tdc_data_ram_0_0_1.REGMODE_A = "NOREG";
    defparam tdc_data_ram_0_0_1.REGMODE_B = "NOREG";
    defparam tdc_data_ram_0_0_1.RESETMODE = "ASYNC";
    defparam tdc_data_ram_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam tdc_data_ram_0_0_1.WRITEMODE_A = "NORMAL";
    defparam tdc_data_ram_0_0_1.WRITEMODE_B = "NORMAL";
    defparam tdc_data_ram_0_0_1.CSDECODE_A = "0b000";
    defparam tdc_data_ram_0_0_1.CSDECODE_B = "0b000";
    defparam tdc_data_ram_0_0_1.GSR = "ENABLED";
    defparam tdc_data_ram_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_0_1.INIT_DATA = "STATIC";
    DP16KD tdc_data_ram_0_1_0 (.DIA0(Data[9]), .DIA1(Data[10]), .DIA2(Data[11]), 
           .DIA3(Data[12]), .DIA4(Data[13]), .DIA5(Data[14]), .DIA6(Data[15]), 
           .DIA7(GND_net), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(WrAddress[0]), .ADA4(WrAddress[1]), 
           .ADA5(WrAddress[2]), .ADA6(WrAddress[3]), .ADA7(WrAddress[4]), 
           .ADA8(WrAddress[5]), .ADA9(WrAddress[6]), .ADA10(WrAddress[7]), 
           .ADA11(WrAddress[8]), .ADA12(WrAddress[9]), .ADA13(WrAddress[10]), 
           .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(Reset), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(GND_net), .ADB3(RdAddress[0]), .ADB4(RdAddress[1]), .ADB5(RdAddress[2]), 
           .ADB6(RdAddress[3]), .ADB7(RdAddress[4]), .ADB8(RdAddress[5]), 
           .ADB9(RdAddress[6]), .ADB10(RdAddress[7]), .ADB11(RdAddress[8]), 
           .ADB12(RdAddress[9]), .ADB13(RdAddress[10]), .CEB(RdClockEn), 
           .OCEB(RdClockEn), .CLKB(RdClock), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(Reset), .DOB0(Q[9]), 
           .DOB1(Q[10]), .DOB2(Q[11]), .DOB3(Q[12]), .DOB4(Q[13]), .DOB5(Q[14]), 
           .DOB6(Q[15])) /* synthesis MEM_LPC_FILE="tdc_data_ram.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;
    defparam tdc_data_ram_0_1_0.DATA_WIDTH_A = 9;
    defparam tdc_data_ram_0_1_0.DATA_WIDTH_B = 9;
    defparam tdc_data_ram_0_1_0.REGMODE_A = "NOREG";
    defparam tdc_data_ram_0_1_0.REGMODE_B = "NOREG";
    defparam tdc_data_ram_0_1_0.RESETMODE = "ASYNC";
    defparam tdc_data_ram_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam tdc_data_ram_0_1_0.WRITEMODE_A = "NORMAL";
    defparam tdc_data_ram_0_1_0.WRITEMODE_B = "NORMAL";
    defparam tdc_data_ram_0_1_0.CSDECODE_A = "0b000";
    defparam tdc_data_ram_0_1_0.CSDECODE_B = "0b000";
    defparam tdc_data_ram_0_1_0.GSR = "ENABLED";
    defparam tdc_data_ram_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam tdc_data_ram_0_1_0.INIT_DATA = "STATIC";
    VHI i13 (.Z(VCC_net));
    GSR GSR_INST (.GSR(VCC_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i4 (.Z(GND_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

